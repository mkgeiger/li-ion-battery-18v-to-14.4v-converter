*****************************************************************************
* DSEI60-06A MACROMODEL *****************************************************
* REV N/A *******************************************************************
*****************************************************************************
*                   ANODE
*                   |  CATHODE
*                   |  |
.SUBCKT  DSEI60-06A 1  2
D1  1  2  DMOD1
.MODEL DMOD1 D (IS=148.21E-6 N=1.8882 RS=3.0622E-3 IKF=811.78E-9 CJO=1.0000E-12 M=.3333 VJ=.75 ISR=406.73E-9 NR=4.9950 BV=600.05 IBV=1.2932E-3 TT=26.602E-9 Vpk=600 Iave=60A mfg=IXYS type=silicon Vpk=600.0V Iave=60.0A)
.ENDS
